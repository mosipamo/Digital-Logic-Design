`timescale 1ns/1ns

module tb_Q7();
    reg [14:0] a = 15'b0;
    wire [3:0] y;

    Q7 u0 (.a(a), .y(y));

    initial begin
	#200
	a[0] = 1;
	#200
	a[1] = 1;
	#200
	a[2] = 1;
	#200
	a[3] = 1;
	#200
	a[4] = 1;
	#200
	a[5] = 1;
	#200
	a[6] = 1;
	#200
	a[7] = 1;
	#200
	a[8] = 1;
	#200
	a[9] = 1;
	#200
	a[10] = 1;
	#200
	a[11] = 1;
	#200
	a[12] = 1;
	#200
	a[13] = 1;
	#200
	a[14] = 1;

	#200			
	a[0] = 0;
	#200
	a[1] = 0;
	#200
	a[2] = 0;
	#200
	a[3] = 0;
	#200
	a[4] = 0;
	#200
	a[5] = 0;
	#200
	a[6] = 0;
	#200
	a[7] = 0;
	#200
	a[8] = 0;
	#200
	a[9] = 0;
	#200
	a[10] = 0;
	#200
	a[11] = 0;
	#200
	a[12] = 0;
	#200
	a[13] = 0;
	#200
	a[14] = 0;
	#200 $stop;
    end
endmodule

